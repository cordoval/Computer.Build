signal22 = '0'